module mem_inst(	
	input clk,
	input  [9:0] addres,
	output [31:0] data_out);
	
  
	reg [31:0] mem [0:1023];
	
		
	always@(*)
		begin
			
		end
	
	assign data_out = mem[addres];
	
endmodule 




/*
j test

			mem[2]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[3]  <=  32'b0000_0100_0000_1000_0000_0000_0111_1000;//li r2 30
			mem[5]  <=  32'b0000_1000_0000_1000_0000_0000_0000_0000;//j 8
			mem[6]  <=  32'b0000_0100_0000_0100_0000_0001_0000_0000;//li r1 64
			mem[8]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//add out r1 r2
	
jr test

			mem[2]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[3]  <=  32'b0000_0100_0000_1000_0000_0000_0010_0100;//li r2 9
			mem[5]  <=  32'b0000_0000_1000_0000_0000_0000_1000_0000;//jr r2
			mem[6]  <=  32'b0000_0100_0000_0100_0000_0001_0000_0000;//li r1 64
			mem[9]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//add out r1 r2
			
jal test

			mem[2]  <=  32'b0000_0100_0000_0100_0000_0000_0100_1000;//li r1 18
			mem[3]  <=  32'b0000_0100_0000_1000_0000_0000_0010_0100;//li r2 9
			mem[5]  <=  32'b0000_1100_0000_1001_0000_0000_0000_0000;//jal 9
			mem[6]  <=  32'b0000_0100_0000_0100_0000_0001_0000_0000;//li r1 64
			mem[9]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//add out r1 r2
			
branch equal test 

			mem[2]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[3]  <=  32'b0000_0100_0000_1000_0000_0000_0111_1000;//li r2 31
			mem[5]  <=  32'b0001_0000_0100_1000_0000_0000_0000_1000;//beq r1 r2 2
			mem[6]  <=  32'b0000_0100_0000_0100_0000_0001_0000_0000;//li r1 64
			mem[8]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//add out r1 r2
			
branch not equal test

			mem[2]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[3]  <=  32'b0000_0100_0000_1000_0000_0000_0111_1100;//li r2 31
			mem[5]  <=  32'b0001_0100_0100_1000_0000_0000_0000_1000;//bne r1 r2 2
			mem[6]  <=  32'b0000_0100_0000_0100_0000_0001_0000_0000;//li r1 64
			mem[8]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//add out r1 r2
sub test

			mem[0]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0010_1100;//li r2 31
			mem[5]  <=  32'b0000_0000_0100_1011_1100_0010_0000_0000;//sub out r1 r2
			
addi test

			mem[0]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0010_1100;//li r2 
			mem[5]  <=  32'b0010_0000_0111_1100_0000_0010_0010_0000;//addi out r1 
			
slti test

			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0101_1000;//li r2 22
			mem[3]  <=  32'b0010_1000_1011_1100_0000_0000_0101_1100;//slti out r2 23
			
slt test

			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0101_1000;//li r2 22
			mem[3]  <=  32'b0000_0000_1000_0111_1100_0010_1010_0000;//slt out s2 s1
			
and + or + sll test

			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0111_0000;//li r1 
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0101_1000;//li r2 
			mem[3]  <=  32'b0000_0000_1000_0100_1100_0010_0100_0000;//and r3 r1 r2
			mem[4]  <=  32'b0000_0000_1000_0111_1100_0010_0101_0000;//or out r1 r2
			mem[5]  <=  32'b0000_0000_0011_1111_1100_1000_0000_0000;//sll out out 2

andi + ori + srl test

			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0111_0000;//li r1 
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0101_1000;//li r2 
			mem[3]  <=  32'b0011_0000_0100_1100_0000_0000_0101_1000;//andi r3 r1 22
			mem[4]  <=  32'b0011_0111_1111_1100_0000_0010_0101_0000;//ori out r1 148
			mem[5]  <=  32'b0000_0000_0011_1111_1100_1000_0010_0000;//srl out out 2
			

SPECIAL TEST-1

			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0111_1000;//li r1 30
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0101_1000;//li r2 22
			mem[3]  <=  32'b1000_1100_0011_1100_0000_0000_0000_1000;//lw out m0(2)
			mem[6]  <=  32'b1010_1100_0000_0100_0000_0000_0000_1000;//sw r1 m0(2)
			mem[8]  <=  32'b1000_1100_0011_1100_0000_0000_0000_1000;//lw out m0(2)
			
SPECIAL TEST-2 
			
			mem[1]  <=  32'b0000_0100_0000_0100_0000_0000_0101_1000;//li r1 22
			mem[2]  <=  32'b0000_0100_0000_1000_0000_0000_0011_1100;//li r2 15
			mem[3]  <=  32'b1000_1100_0000_1000_0000_0000_0001_0000;//sw r2  m0(4)
			mem[6]  <=  32'b1010_1100_0000_0100_0000_0000_0000_1000;//sw r1  m0(2)
			mem[8]  <=  32'b1000_1100_0000_1100_0000_0000_0001_0000;//lw r3  m0(4)
			mem[11] <=  32'b1000_1100_0011_1100_0000_0000_0000_1000;//lw out m0(2)
			mem[8]  <=  32'b0000_0000_1111_1111_1100_0010_0000_0000;//add out out r3
			
*/



