module c_r(
	input s,
	output out);
	
	or or1(out , s , 0);
	
endmodule 