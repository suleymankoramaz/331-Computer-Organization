module and32(
				input  [31:0] a,
				input  [31:0] b,
				output [31:0] out);

	and and1( out[0]  , a[0]  , b[0]);
	and and2( out[1]  , a[1]  , b[1]);
	and and3( out[2]  , a[2]  , b[2]);
	and and4( out[3]  , a[3]  , b[3]);
	and and5( out[4]  , a[4]  , b[4]);
	and and6( out[5]  , a[5]  , b[5]);
	and and7( out[6]  , a[6]  , b[6]);
	and and8( out[7]  , a[7]  , b[7]);
	and and9( out[8]  , a[8]  , b[8]);
	and and10(out[9]  , a[9]  , b[9]);
	and and11(out[10] , a[10] , b[10]);
	and and12(out[11] , a[11] , b[11]);
	and and13(out[12] , a[12] , b[12]);
	and and14(out[13] , a[13] , b[13]);
	and and15(out[14] , a[14] , b[14]);
	and and16(out[15] , a[15] , b[15]);
	and and17(out[16] , a[16] , b[16]);
	and and18(out[17] , a[17] , b[17]);
	and and19(out[18] , a[18] , b[18]);
	and and20(out[19] , a[19] , b[19]);
	and and21(out[20] , a[20] , b[20]);
	and and22(out[21] , a[21] , b[21]);
	and and23(out[22] , a[22] , b[22]);
	and and24(out[23] , a[23] , b[23]);
	and and25(out[24] , a[24] , b[24]);
	and and26(out[25] , a[25] , b[25]);
	and and27(out[26] , a[26] , b[26]);
	and and28(out[27] , a[27] , b[27]);
	and and29(out[28] , a[28] , b[28]);
	and and30(out[29] , a[29] , b[29]);
	and and31(out[30] , a[30] , b[30]);
	and and32(out[31] , a[31] , b[31]);
endmodule